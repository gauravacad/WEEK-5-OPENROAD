module gcd (clk,
    req_rdy,
    req_val,
    reset,
    resp_rdy,
    resp_val,
    req_msg,
    resp_msg);
 input clk;
 output req_rdy;
 input req_val;
 input reset;
 input resp_rdy;
 output resp_val;
 input [31:0] req_msg;
 output [15:0] resp_msg;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _167_;
 wire _168_;
 wire _172_;
 wire _174_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _190_;
 wire _191_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire net2;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire net1;
 wire _235_;
 wire _236_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire \ctrl.state.out[1] ;
 wire \ctrl.state.out[2] ;
 wire \dpath.a_lt_b$in0[0] ;
 wire \dpath.a_lt_b$in0[10] ;
 wire \dpath.a_lt_b$in0[11] ;
 wire \dpath.a_lt_b$in0[12] ;
 wire \dpath.a_lt_b$in0[13] ;
 wire \dpath.a_lt_b$in0[14] ;
 wire \dpath.a_lt_b$in0[15] ;
 wire \dpath.a_lt_b$in0[1] ;
 wire \dpath.a_lt_b$in0[2] ;
 wire \dpath.a_lt_b$in0[3] ;
 wire \dpath.a_lt_b$in0[4] ;
 wire \dpath.a_lt_b$in0[5] ;
 wire \dpath.a_lt_b$in0[6] ;
 wire \dpath.a_lt_b$in0[7] ;
 wire \dpath.a_lt_b$in0[8] ;
 wire \dpath.a_lt_b$in0[9] ;
 wire \dpath.a_lt_b$in1[0] ;
 wire \dpath.a_lt_b$in1[10] ;
 wire \dpath.a_lt_b$in1[11] ;
 wire \dpath.a_lt_b$in1[12] ;
 wire \dpath.a_lt_b$in1[13] ;
 wire \dpath.a_lt_b$in1[14] ;
 wire \dpath.a_lt_b$in1[15] ;
 wire \dpath.a_lt_b$in1[1] ;
 wire \dpath.a_lt_b$in1[2] ;
 wire \dpath.a_lt_b$in1[3] ;
 wire \dpath.a_lt_b$in1[4] ;
 wire \dpath.a_lt_b$in1[5] ;
 wire \dpath.a_lt_b$in1[6] ;
 wire \dpath.a_lt_b$in1[7] ;
 wire \dpath.a_lt_b$in1[8] ;
 wire \dpath.a_lt_b$in1[9] ;

 INV_X2 _345_ (.A(\dpath.a_lt_b$in1[1] ),
    .ZN(_036_));
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 NAND2_X1 _347_ (.A1(_036_),
    .A2(\dpath.a_lt_b$in0[1] ),
    .ZN(_038_));
 INV_X1 _348_ (.A(\dpath.a_lt_b$in1[0] ),
    .ZN(_039_));
 NOR2_X1 _349_ (.A1(_039_),
    .A2(\dpath.a_lt_b$in0[0] ),
    .ZN(_040_));
 NOR2_X1 _350_ (.A1(_036_),
    .A2(\dpath.a_lt_b$in0[1] ),
    .ZN(_041_));
 OAI21_X2 _351_ (.A(_038_),
    .B1(_040_),
    .B2(_041_),
    .ZN(_042_));
 INV_X1 _352_ (.A(\dpath.a_lt_b$in1[3] ),
    .ZN(_043_));
 NAND2_X1 _353_ (.A1(_043_),
    .A2(\dpath.a_lt_b$in0[3] ),
    .ZN(_044_));
 INV_X1 _354_ (.A(\dpath.a_lt_b$in0[3] ),
    .ZN(_045_));
 NAND2_X1 _355_ (.A1(_045_),
    .A2(\dpath.a_lt_b$in1[3] ),
    .ZN(_046_));
 NAND2_X1 _356_ (.A1(_044_),
    .A2(_046_),
    .ZN(_047_));
 INV_X2 _357_ (.A(\dpath.a_lt_b$in1[2] ),
    .ZN(_048_));
 NAND2_X2 _358_ (.A1(_048_),
    .A2(\dpath.a_lt_b$in0[2] ),
    .ZN(_049_));
 INV_X1 _359_ (.A(\dpath.a_lt_b$in0[2] ),
    .ZN(_050_));
 NAND2_X1 _360_ (.A1(_050_),
    .A2(\dpath.a_lt_b$in1[2] ),
    .ZN(_051_));
 NAND2_X2 _361_ (.A1(_049_),
    .A2(_051_),
    .ZN(_052_));
 NOR2_X2 _362_ (.A1(_047_),
    .A2(_052_),
    .ZN(_053_));
 NAND2_X2 _363_ (.A1(_042_),
    .A2(_053_),
    .ZN(_054_));
 INV_X1 _364_ (.A(_046_),
    .ZN(_055_));
 OAI21_X1 _365_ (.A(_044_),
    .B1(_055_),
    .B2(_049_),
    .ZN(_056_));
 INV_X1 _366_ (.A(_056_),
    .ZN(_057_));
 NAND2_X4 _367_ (.A1(_054_),
    .A2(_057_),
    .ZN(_058_));
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 XNOR2_X2 _369_ (.A(\dpath.a_lt_b$in1[5] ),
    .B(\dpath.a_lt_b$in0[5] ),
    .ZN(_060_));
 XNOR2_X1 _370_ (.A(\dpath.a_lt_b$in1[4] ),
    .B(\dpath.a_lt_b$in0[4] ),
    .ZN(_061_));
 NAND2_X1 _371_ (.A1(_060_),
    .A2(_061_),
    .ZN(_062_));
 XNOR2_X2 _372_ (.A(\dpath.a_lt_b$in1[7] ),
    .B(\dpath.a_lt_b$in0[7] ),
    .ZN(_063_));
 XNOR2_X2 _373_ (.A(\dpath.a_lt_b$in1[6] ),
    .B(\dpath.a_lt_b$in0[6] ),
    .ZN(_064_));
 NAND2_X1 _374_ (.A1(_063_),
    .A2(_064_),
    .ZN(_065_));
 NOR2_X1 _375_ (.A1(_062_),
    .A2(_065_),
    .ZN(_066_));
 NAND2_X2 _376_ (.A1(_058_),
    .A2(_066_),
    .ZN(_067_));
 INV_X1 _377_ (.A(\dpath.a_lt_b$in1[4] ),
    .ZN(_068_));
 NAND2_X1 _378_ (.A1(_068_),
    .A2(\dpath.a_lt_b$in0[4] ),
    .ZN(_069_));
 INV_X1 _379_ (.A(\dpath.a_lt_b$in0[5] ),
    .ZN(_070_));
 OAI21_X2 _380_ (.A(_069_),
    .B1(\dpath.a_lt_b$in1[5] ),
    .B2(_070_),
    .ZN(_071_));
 INV_X1 _381_ (.A(\dpath.a_lt_b$in1[5] ),
    .ZN(_072_));
 NOR2_X2 _382_ (.A1(_072_),
    .A2(\dpath.a_lt_b$in0[5] ),
    .ZN(_073_));
 INV_X1 _383_ (.A(_073_),
    .ZN(_074_));
 NAND2_X1 _384_ (.A1(_071_),
    .A2(_074_),
    .ZN(_075_));
 NOR2_X1 _385_ (.A1(_075_),
    .A2(_065_),
    .ZN(_076_));
 INV_X1 _386_ (.A(\dpath.a_lt_b$in1[7] ),
    .ZN(_077_));
 NAND2_X1 _387_ (.A1(_077_),
    .A2(\dpath.a_lt_b$in0[7] ),
    .ZN(_078_));
 INV_X2 _388_ (.A(_063_),
    .ZN(_079_));
 INV_X1 _389_ (.A(\dpath.a_lt_b$in1[6] ),
    .ZN(_080_));
 NAND2_X1 _390_ (.A1(_080_),
    .A2(\dpath.a_lt_b$in0[6] ),
    .ZN(_081_));
 OAI21_X1 _391_ (.A(_078_),
    .B1(_079_),
    .B2(_081_),
    .ZN(_082_));
 NOR2_X2 _392_ (.A1(_076_),
    .A2(_082_),
    .ZN(_083_));
 NAND2_X4 _393_ (.A1(_067_),
    .A2(_083_),
    .ZN(_084_));
 INV_X2 _394_ (.A(\dpath.a_lt_b$in1[11] ),
    .ZN(_085_));
 XNOR2_X2 _395_ (.A(_085_),
    .B(\dpath.a_lt_b$in0[11] ),
    .ZN(_086_));
 INV_X2 _396_ (.A(\dpath.a_lt_b$in1[10] ),
    .ZN(_087_));
 XNOR2_X1 _397_ (.A(_087_),
    .B(\dpath.a_lt_b$in0[10] ),
    .ZN(_088_));
 NOR2_X2 _398_ (.A1(_086_),
    .A2(_088_),
    .ZN(_089_));
 XNOR2_X2 _399_ (.A(\dpath.a_lt_b$in1[9] ),
    .B(\dpath.a_lt_b$in0[9] ),
    .ZN(_090_));
 XNOR2_X2 _400_ (.A(\dpath.a_lt_b$in1[8] ),
    .B(\dpath.a_lt_b$in0[8] ),
    .ZN(_091_));
 NAND2_X1 _401_ (.A1(_090_),
    .A2(_091_),
    .ZN(_092_));
 INV_X1 _402_ (.A(_092_),
    .ZN(_093_));
 AND2_X1 _403_ (.A1(_089_),
    .A2(_093_),
    .ZN(_094_));
 NAND2_X2 _404_ (.A1(_084_),
    .A2(_094_),
    .ZN(_095_));
 NAND2_X1 _405_ (.A1(_085_),
    .A2(\dpath.a_lt_b$in0[11] ),
    .ZN(_096_));
 NAND2_X1 _406_ (.A1(_087_),
    .A2(\dpath.a_lt_b$in0[10] ),
    .ZN(_097_));
 OAI21_X1 _407_ (.A(_096_),
    .B1(_086_),
    .B2(_097_),
    .ZN(_098_));
 INV_X1 _408_ (.A(\dpath.a_lt_b$in0[9] ),
    .ZN(_099_));
 NOR2_X1 _409_ (.A1(_099_),
    .A2(\dpath.a_lt_b$in1[9] ),
    .ZN(_100_));
 INV_X1 _410_ (.A(\dpath.a_lt_b$in1[8] ),
    .ZN(_101_));
 AND2_X1 _411_ (.A1(_101_),
    .A2(\dpath.a_lt_b$in0[8] ),
    .ZN(_102_));
 AOI21_X2 _412_ (.A(_100_),
    .B1(_090_),
    .B2(_102_),
    .ZN(_103_));
 INV_X1 _413_ (.A(_103_),
    .ZN(_104_));
 AOI21_X2 _414_ (.A(_098_),
    .B1(_104_),
    .B2(_089_),
    .ZN(_105_));
 NAND2_X4 _415_ (.A1(_095_),
    .A2(_105_),
    .ZN(_106_));
 XNOR2_X2 _416_ (.A(\dpath.a_lt_b$in1[12] ),
    .B(\dpath.a_lt_b$in0[12] ),
    .ZN(_107_));
 INV_X1 _417_ (.A(_107_),
    .ZN(_108_));
 INV_X2 _418_ (.A(\dpath.a_lt_b$in1[13] ),
    .ZN(_109_));
 XNOR2_X2 _419_ (.A(_109_),
    .B(\dpath.a_lt_b$in0[13] ),
    .ZN(_110_));
 NOR2_X2 _420_ (.A1(_108_),
    .A2(_110_),
    .ZN(_111_));
 NAND2_X2 _421_ (.A1(_106_),
    .A2(_111_),
    .ZN(_112_));
 NAND2_X1 _422_ (.A1(_109_),
    .A2(\dpath.a_lt_b$in0[13] ),
    .ZN(_113_));
 INV_X1 _423_ (.A(\dpath.a_lt_b$in1[12] ),
    .ZN(_114_));
 NAND2_X1 _424_ (.A1(_114_),
    .A2(\dpath.a_lt_b$in0[12] ),
    .ZN(_115_));
 OAI21_X1 _425_ (.A(_113_),
    .B1(_110_),
    .B2(_115_),
    .ZN(_116_));
 INV_X1 _426_ (.A(_116_),
    .ZN(_117_));
 NAND2_X2 _427_ (.A1(_112_),
    .A2(_117_),
    .ZN(_118_));
 INV_X1 _428_ (.A(\dpath.a_lt_b$in1[14] ),
    .ZN(_119_));
 XNOR2_X1 _429_ (.A(_119_),
    .B(\dpath.a_lt_b$in0[14] ),
    .ZN(_120_));
 INV_X1 _430_ (.A(_120_),
    .ZN(_121_));
 NAND2_X2 _431_ (.A1(_118_),
    .A2(_121_),
    .ZN(_122_));
 NAND2_X1 _432_ (.A1(_119_),
    .A2(\dpath.a_lt_b$in0[14] ),
    .ZN(_123_));
 NAND2_X1 _433_ (.A1(_122_),
    .A2(_123_),
    .ZN(_124_));
 INV_X2 _434_ (.A(\dpath.a_lt_b$in1[15] ),
    .ZN(_125_));
 XNOR2_X1 _435_ (.A(_125_),
    .B(\dpath.a_lt_b$in0[15] ),
    .ZN(_126_));
 INV_X1 _436_ (.A(_126_),
    .ZN(_127_));
 NAND2_X1 _437_ (.A1(_124_),
    .A2(_127_),
    .ZN(_128_));
 NAND3_X1 _438_ (.A1(_122_),
    .A2(_123_),
    .A3(_126_),
    .ZN(_129_));
 AND2_X1 _439_ (.A1(_128_),
    .A2(_129_),
    .ZN(resp_msg[15]));
 XNOR2_X1 _440_ (.A(\dpath.a_lt_b$in1[1] ),
    .B(\dpath.a_lt_b$in0[1] ),
    .ZN(_130_));
 INV_X1 _441_ (.A(_040_),
    .ZN(_131_));
 XNOR2_X1 _442_ (.A(_130_),
    .B(_131_),
    .ZN(_132_));
 INV_X1 _443_ (.A(_132_),
    .ZN(resp_msg[1]));
 INV_X1 _444_ (.A(_052_),
    .ZN(_133_));
 XNOR2_X1 _445_ (.A(_042_),
    .B(_133_),
    .ZN(_134_));
 INV_X1 _446_ (.A(_134_),
    .ZN(resp_msg[2]));
 NAND2_X1 _447_ (.A1(_042_),
    .A2(_133_),
    .ZN(_135_));
 NAND2_X1 _448_ (.A1(_135_),
    .A2(_049_),
    .ZN(_136_));
 XNOR2_X1 _449_ (.A(_136_),
    .B(_047_),
    .ZN(resp_msg[3]));
 XNOR2_X1 _450_ (.A(_058_),
    .B(_061_),
    .ZN(_137_));
 INV_X1 _451_ (.A(_137_),
    .ZN(resp_msg[4]));
 NAND2_X1 _452_ (.A1(_058_),
    .A2(_061_),
    .ZN(_138_));
 NAND2_X1 _453_ (.A1(_138_),
    .A2(_069_),
    .ZN(_139_));
 XOR2_X1 _454_ (.A(_139_),
    .B(_060_),
    .Z(resp_msg[5]));
 INV_X1 _455_ (.A(_071_),
    .ZN(_140_));
 AOI21_X2 _456_ (.A(_073_),
    .B1(_138_),
    .B2(_140_),
    .ZN(_141_));
 XNOR2_X1 _457_ (.A(_141_),
    .B(_064_),
    .ZN(_142_));
 INV_X1 _458_ (.A(_142_),
    .ZN(resp_msg[6]));
 NAND2_X1 _459_ (.A1(_141_),
    .A2(_064_),
    .ZN(_143_));
 NAND2_X1 _460_ (.A1(_143_),
    .A2(_081_),
    .ZN(_144_));
 XNOR2_X1 _461_ (.A(_144_),
    .B(_079_),
    .ZN(resp_msg[7]));
 XNOR2_X1 _462_ (.A(_084_),
    .B(_091_),
    .ZN(_145_));
 INV_X1 _463_ (.A(_145_),
    .ZN(resp_msg[8]));
 AOI21_X1 _464_ (.A(_102_),
    .B1(_084_),
    .B2(_091_),
    .ZN(_146_));
 XNOR2_X1 _465_ (.A(_146_),
    .B(_090_),
    .ZN(resp_msg[9]));
 NAND2_X1 _466_ (.A1(_084_),
    .A2(_093_),
    .ZN(_147_));
 NAND2_X2 _467_ (.A1(_147_),
    .A2(_103_),
    .ZN(_148_));
 INV_X1 _468_ (.A(_088_),
    .ZN(_149_));
 XNOR2_X1 _469_ (.A(_148_),
    .B(_149_),
    .ZN(_150_));
 INV_X1 _470_ (.A(_150_),
    .ZN(resp_msg[10]));
 NAND2_X2 _471_ (.A1(_148_),
    .A2(_149_),
    .ZN(_151_));
 NAND2_X2 _472_ (.A1(_151_),
    .A2(_097_),
    .ZN(_152_));
 XNOR2_X2 _473_ (.A(_152_),
    .B(_086_),
    .ZN(resp_msg[11]));
 XNOR2_X1 _474_ (.A(_106_),
    .B(_107_),
    .ZN(_153_));
 INV_X1 _475_ (.A(_153_),
    .ZN(resp_msg[12]));
 NAND2_X2 _476_ (.A1(_106_),
    .A2(_107_),
    .ZN(_154_));
 NAND2_X2 _477_ (.A1(_154_),
    .A2(_115_),
    .ZN(_155_));
 XNOR2_X2 _478_ (.A(_155_),
    .B(_110_),
    .ZN(resp_msg[13]));
 XNOR2_X1 _479_ (.A(_118_),
    .B(_121_),
    .ZN(_156_));
 INV_X1 _480_ (.A(_156_),
    .ZN(resp_msg[14]));
 XNOR2_X1 _481_ (.A(_039_),
    .B(\dpath.a_lt_b$in0[0] ),
    .ZN(resp_msg[0]));
 NAND4_X1 _482_ (.A1(_119_),
    .A2(_125_),
    .A3(_039_),
    .A4(_036_),
    .ZN(_157_));
 NAND3_X1 _483_ (.A1(_087_),
    .A2(_085_),
    .A3(_114_),
    .ZN(_158_));
 NOR3_X1 _484_ (.A1(_157_),
    .A2(\dpath.a_lt_b$in1[13] ),
    .A3(_158_),
    .ZN(_159_));
 INV_X1 _485_ (.A(\dpath.a_lt_b$in1[9] ),
    .ZN(_160_));
 NAND4_X1 _486_ (.A1(_080_),
    .A2(_077_),
    .A3(_101_),
    .A4(_160_),
    .ZN(_161_));
 NAND4_X1 _487_ (.A1(_048_),
    .A2(_043_),
    .A3(_068_),
    .A4(_072_),
    .ZN(_162_));
 NOR2_X1 _488_ (.A1(_161_),
    .A2(_162_),
    .ZN(_163_));
 NAND2_X1 _489_ (.A1(_159_),
    .A2(_163_),
    .ZN(_164_));
 INV_X1 _490_ (.A(_164_),
    .ZN(_165_));
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 INV_X1 _492_ (.A(\ctrl.state.out[2] ),
    .ZN(_167_));
 OR2_X1 _493_ (.A1(_167_),
    .A2(reset),
    .ZN(_168_));
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 NAND2_X1 _497_ (.A1(req_rdy),
    .A2(req_val),
    .ZN(_172_));
 OAI22_X1 _498_ (.A1(_165_),
    .A2(_168_),
    .B1(reset),
    .B2(_172_),
    .ZN(_002_));
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 AND3_X1 _500_ (.A1(_167_),
    .A2(_003_),
    .A3(\ctrl.state.out[1] ),
    .ZN(resp_val));
 AOI21_X1 _501_ (.A(reset),
    .B1(resp_val),
    .B2(resp_rdy),
    .ZN(_174_));
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 INV_X1 _503_ (.A(req_rdy),
    .ZN(_176_));
 OAI21_X1 _504_ (.A(_174_),
    .B1(_176_),
    .B2(req_val),
    .ZN(_000_));
 NAND2_X1 _505_ (.A1(_174_),
    .A2(\ctrl.state.out[1] ),
    .ZN(_177_));
 OAI21_X1 _506_ (.A(_177_),
    .B1(_164_),
    .B2(_168_),
    .ZN(_001_));
 NAND2_X1 _507_ (.A1(_125_),
    .A2(\dpath.a_lt_b$in0[15] ),
    .ZN(_178_));
 OAI21_X1 _508_ (.A(_178_),
    .B1(_126_),
    .B2(_123_),
    .ZN(_179_));
 NOR2_X2 _509_ (.A1(_120_),
    .A2(_126_),
    .ZN(_180_));
 AOI21_X1 _510_ (.A(_179_),
    .B1(_116_),
    .B2(_180_),
    .ZN(_181_));
 NAND2_X1 _511_ (.A1(_111_),
    .A2(_180_),
    .ZN(_182_));
 OAI21_X1 _512_ (.A(_181_),
    .B1(_105_),
    .B2(_182_),
    .ZN(_183_));
 INV_X2 _513_ (.A(_183_),
    .ZN(_184_));
 INV_X1 _514_ (.A(_182_),
    .ZN(_185_));
 NAND3_X4 _515_ (.A1(_084_),
    .A2(_094_),
    .A3(_185_),
    .ZN(_186_));
 NAND3_X1 _516_ (.A1(_184_),
    .A2(_186_),
    .A3(\ctrl.state.out[2] ),
    .ZN(_187_));
 NAND2_X2 _517_ (.A1(_187_),
    .A2(_003_),
    .ZN(_188_));
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 MUX2_X1 _519_ (.A(\dpath.a_lt_b$in0[0] ),
    .B(req_msg[0]),
    .S(net2),
    .Z(_190_));
 NAND2_X1 _520_ (.A1(_188_),
    .A2(_190_),
    .ZN(_191_));
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 OAI21_X1 _522_ (.A(_191_),
    .B1(_039_),
    .B2(_188_),
    .ZN(_004_));
 MUX2_X1 _523_ (.A(\dpath.a_lt_b$in0[1] ),
    .B(req_msg[1]),
    .S(net2),
    .Z(_193_));
 NAND2_X1 _524_ (.A1(_188_),
    .A2(_193_),
    .ZN(_194_));
 OAI21_X1 _525_ (.A(_194_),
    .B1(_036_),
    .B2(_188_),
    .ZN(_005_));
 NAND2_X1 _526_ (.A1(req_rdy),
    .A2(req_msg[2]),
    .ZN(_195_));
 OAI21_X1 _527_ (.A(_195_),
    .B1(req_rdy),
    .B2(_050_),
    .ZN(_196_));
 NAND2_X1 _528_ (.A1(_188_),
    .A2(_196_),
    .ZN(_197_));
 OAI21_X1 _529_ (.A(_197_),
    .B1(_048_),
    .B2(_188_),
    .ZN(_006_));
 NAND2_X1 _530_ (.A1(req_rdy),
    .A2(req_msg[3]),
    .ZN(_198_));
 OAI21_X1 _531_ (.A(_198_),
    .B1(req_rdy),
    .B2(_045_),
    .ZN(_199_));
 NAND2_X1 _532_ (.A1(_188_),
    .A2(_199_),
    .ZN(_200_));
 OAI21_X1 _533_ (.A(_200_),
    .B1(_043_),
    .B2(_188_),
    .ZN(_007_));
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 MUX2_X1 _536_ (.A(\dpath.a_lt_b$in0[4] ),
    .B(req_msg[4]),
    .S(req_rdy),
    .Z(_203_));
 NAND2_X1 _537_ (.A1(_188_),
    .A2(_203_),
    .ZN(_204_));
 OAI21_X1 _538_ (.A(_204_),
    .B1(_068_),
    .B2(_188_),
    .ZN(_008_));
 NAND2_X1 _539_ (.A1(req_rdy),
    .A2(req_msg[5]),
    .ZN(_205_));
 OAI21_X1 _540_ (.A(_205_),
    .B1(req_rdy),
    .B2(_070_),
    .ZN(_206_));
 NAND2_X1 _541_ (.A1(_188_),
    .A2(_206_),
    .ZN(_207_));
 OAI21_X1 _542_ (.A(_207_),
    .B1(_072_),
    .B2(_188_),
    .ZN(_009_));
 MUX2_X1 _543_ (.A(\dpath.a_lt_b$in0[6] ),
    .B(req_msg[6]),
    .S(req_rdy),
    .Z(_208_));
 NAND2_X1 _544_ (.A1(_188_),
    .A2(_208_),
    .ZN(_209_));
 OAI21_X1 _545_ (.A(_209_),
    .B1(_080_),
    .B2(_188_),
    .ZN(_010_));
 MUX2_X1 _546_ (.A(\dpath.a_lt_b$in0[7] ),
    .B(req_msg[7]),
    .S(req_rdy),
    .Z(_210_));
 NAND2_X1 _547_ (.A1(_188_),
    .A2(_210_),
    .ZN(_211_));
 OAI21_X1 _548_ (.A(_211_),
    .B1(_077_),
    .B2(_188_),
    .ZN(_011_));
 MUX2_X1 _549_ (.A(\dpath.a_lt_b$in0[8] ),
    .B(req_msg[8]),
    .S(req_rdy),
    .Z(_212_));
 NAND2_X1 _550_ (.A1(_188_),
    .A2(_212_),
    .ZN(_213_));
 OAI21_X1 _551_ (.A(_213_),
    .B1(_101_),
    .B2(_188_),
    .ZN(_012_));
 NAND2_X1 _552_ (.A1(req_rdy),
    .A2(req_msg[9]),
    .ZN(_214_));
 OAI21_X1 _553_ (.A(_214_),
    .B1(req_rdy),
    .B2(_099_),
    .ZN(_215_));
 NAND2_X1 _554_ (.A1(_188_),
    .A2(_215_),
    .ZN(_216_));
 OAI21_X1 _555_ (.A(_216_),
    .B1(_160_),
    .B2(_188_),
    .ZN(_013_));
 MUX2_X1 _556_ (.A(\dpath.a_lt_b$in0[10] ),
    .B(req_msg[10]),
    .S(req_rdy),
    .Z(_217_));
 NAND2_X1 _557_ (.A1(_188_),
    .A2(_217_),
    .ZN(_218_));
 OAI21_X1 _558_ (.A(_218_),
    .B1(_087_),
    .B2(_188_),
    .ZN(_014_));
 MUX2_X1 _559_ (.A(\dpath.a_lt_b$in0[11] ),
    .B(req_msg[11]),
    .S(req_rdy),
    .Z(_219_));
 NAND2_X1 _560_ (.A1(_188_),
    .A2(_219_),
    .ZN(_220_));
 OAI21_X1 _561_ (.A(_220_),
    .B1(_085_),
    .B2(_188_),
    .ZN(_015_));
 MUX2_X1 _562_ (.A(\dpath.a_lt_b$in0[12] ),
    .B(req_msg[12]),
    .S(net2),
    .Z(_221_));
 NAND2_X1 _563_ (.A1(_188_),
    .A2(_221_),
    .ZN(_222_));
 OAI21_X1 _564_ (.A(_222_),
    .B1(_114_),
    .B2(_188_),
    .ZN(_016_));
 MUX2_X1 _565_ (.A(\dpath.a_lt_b$in0[13] ),
    .B(req_msg[13]),
    .S(net2),
    .Z(_223_));
 NAND2_X1 _566_ (.A1(_188_),
    .A2(_223_),
    .ZN(_224_));
 OAI21_X1 _567_ (.A(_224_),
    .B1(_109_),
    .B2(_188_),
    .ZN(_017_));
 MUX2_X1 _568_ (.A(\dpath.a_lt_b$in0[14] ),
    .B(req_msg[14]),
    .S(net2),
    .Z(_225_));
 NAND2_X1 _569_ (.A1(_188_),
    .A2(_225_),
    .ZN(_226_));
 OAI21_X1 _570_ (.A(_226_),
    .B1(_119_),
    .B2(_188_),
    .ZN(_018_));
 MUX2_X1 _571_ (.A(\dpath.a_lt_b$in0[15] ),
    .B(req_msg[15]),
    .S(net2),
    .Z(_227_));
 NAND2_X1 _572_ (.A1(_188_),
    .A2(_227_),
    .ZN(_228_));
 OAI21_X1 _573_ (.A(_228_),
    .B1(_125_),
    .B2(_188_),
    .ZN(_019_));
 NAND2_X4 _574_ (.A1(_184_),
    .A2(_186_),
    .ZN(_229_));
 NAND3_X4 _575_ (.A1(_229_),
    .A2(\ctrl.state.out[2] ),
    .A3(_003_),
    .ZN(_230_));
 INV_X8 _576_ (.A(_230_),
    .ZN(_231_));
 NAND2_X1 _577_ (.A1(_231_),
    .A2(resp_msg[0]),
    .ZN(_232_));
 NAND4_X4 _578_ (.A1(_184_),
    .A2(_186_),
    .A3(\ctrl.state.out[2] ),
    .A4(_003_),
    .ZN(_233_));
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 OAI21_X1 _580_ (.A(_232_),
    .B1(_233_),
    .B2(_039_),
    .ZN(_235_));
 NOR2_X2 _581_ (.A1(_167_),
    .A2(req_rdy),
    .ZN(_236_));
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 NAND2_X1 _583_ (.A1(_235_),
    .A2(_236_),
    .ZN(_238_));
 NAND2_X1 _584_ (.A1(net2),
    .A2(req_msg[16]),
    .ZN(_239_));
 NOR2_X1 _585_ (.A1(\ctrl.state.out[2] ),
    .A2(req_rdy),
    .ZN(_240_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 NAND2_X1 _587_ (.A1(net1),
    .A2(\dpath.a_lt_b$in0[0] ),
    .ZN(_242_));
 NAND3_X1 _588_ (.A1(_238_),
    .A2(_239_),
    .A3(_242_),
    .ZN(_020_));
 OAI22_X1 _589_ (.A1(_233_),
    .A2(_036_),
    .B1(_230_),
    .B2(_132_),
    .ZN(_243_));
 NAND2_X1 _590_ (.A1(_243_),
    .A2(_236_),
    .ZN(_244_));
 NAND2_X1 _591_ (.A1(net2),
    .A2(req_msg[17]),
    .ZN(_245_));
 NAND2_X1 _592_ (.A1(net1),
    .A2(\dpath.a_lt_b$in0[1] ),
    .ZN(_246_));
 NAND3_X1 _593_ (.A1(_244_),
    .A2(_245_),
    .A3(_246_),
    .ZN(_021_));
 OAI22_X1 _594_ (.A1(_233_),
    .A2(_048_),
    .B1(_230_),
    .B2(_134_),
    .ZN(_247_));
 NAND2_X1 _595_ (.A1(_247_),
    .A2(_236_),
    .ZN(_248_));
 NAND2_X1 _596_ (.A1(req_msg[18]),
    .A2(req_rdy),
    .ZN(_249_));
 NAND2_X1 _597_ (.A1(net1),
    .A2(\dpath.a_lt_b$in0[2] ),
    .ZN(_250_));
 NAND3_X1 _598_ (.A1(_248_),
    .A2(_249_),
    .A3(_250_),
    .ZN(_022_));
 NAND2_X1 _599_ (.A1(_231_),
    .A2(resp_msg[3]),
    .ZN(_251_));
 OAI21_X1 _600_ (.A(_251_),
    .B1(_233_),
    .B2(_043_),
    .ZN(_252_));
 NAND2_X1 _601_ (.A1(_252_),
    .A2(_236_),
    .ZN(_253_));
 NAND2_X1 _602_ (.A1(req_msg[19]),
    .A2(req_rdy),
    .ZN(_254_));
 NAND2_X1 _603_ (.A1(net1),
    .A2(\dpath.a_lt_b$in0[3] ),
    .ZN(_255_));
 NAND3_X1 _604_ (.A1(_253_),
    .A2(_254_),
    .A3(_255_),
    .ZN(_023_));
 OAI22_X1 _605_ (.A1(_233_),
    .A2(_068_),
    .B1(_230_),
    .B2(_137_),
    .ZN(_256_));
 NAND2_X1 _606_ (.A1(_256_),
    .A2(_236_),
    .ZN(_257_));
 NAND2_X1 _607_ (.A1(req_msg[20]),
    .A2(req_rdy),
    .ZN(_258_));
 NAND2_X1 _608_ (.A1(net1),
    .A2(\dpath.a_lt_b$in0[4] ),
    .ZN(_259_));
 NAND3_X1 _609_ (.A1(_257_),
    .A2(_258_),
    .A3(_259_),
    .ZN(_024_));
 NAND2_X1 _610_ (.A1(_231_),
    .A2(resp_msg[5]),
    .ZN(_260_));
 OAI21_X1 _611_ (.A(_260_),
    .B1(_233_),
    .B2(_072_),
    .ZN(_261_));
 NAND2_X1 _612_ (.A1(_261_),
    .A2(_236_),
    .ZN(_262_));
 NAND2_X1 _613_ (.A1(req_msg[21]),
    .A2(req_rdy),
    .ZN(_263_));
 NAND2_X1 _614_ (.A1(net1),
    .A2(\dpath.a_lt_b$in0[5] ),
    .ZN(_264_));
 NAND3_X1 _615_ (.A1(_262_),
    .A2(_263_),
    .A3(_264_),
    .ZN(_025_));
 OAI22_X1 _616_ (.A1(_233_),
    .A2(_080_),
    .B1(_230_),
    .B2(_142_),
    .ZN(_265_));
 NAND2_X1 _617_ (.A1(_265_),
    .A2(_236_),
    .ZN(_266_));
 NAND2_X1 _618_ (.A1(req_msg[22]),
    .A2(req_rdy),
    .ZN(_267_));
 NAND2_X1 _619_ (.A1(net1),
    .A2(\dpath.a_lt_b$in0[6] ),
    .ZN(_268_));
 NAND3_X1 _620_ (.A1(_266_),
    .A2(_267_),
    .A3(_268_),
    .ZN(_026_));
 NAND2_X1 _621_ (.A1(resp_msg[7]),
    .A2(_231_),
    .ZN(_269_));
 OAI21_X1 _622_ (.A(_269_),
    .B1(_077_),
    .B2(_233_),
    .ZN(_270_));
 NAND2_X1 _623_ (.A1(_270_),
    .A2(_236_),
    .ZN(_271_));
 NAND2_X1 _624_ (.A1(req_msg[23]),
    .A2(req_rdy),
    .ZN(_272_));
 NAND2_X1 _625_ (.A1(net1),
    .A2(\dpath.a_lt_b$in0[7] ),
    .ZN(_273_));
 NAND3_X1 _626_ (.A1(_271_),
    .A2(_272_),
    .A3(_273_),
    .ZN(_027_));
 OAI22_X1 _627_ (.A1(_233_),
    .A2(_101_),
    .B1(_230_),
    .B2(_145_),
    .ZN(_274_));
 NAND2_X1 _628_ (.A1(_274_),
    .A2(_236_),
    .ZN(_275_));
 NAND2_X1 _629_ (.A1(req_msg[24]),
    .A2(req_rdy),
    .ZN(_276_));
 NAND2_X1 _630_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[8] ),
    .ZN(_277_));
 NAND3_X1 _631_ (.A1(_275_),
    .A2(_276_),
    .A3(_277_),
    .ZN(_028_));
 NAND2_X1 _632_ (.A1(_231_),
    .A2(resp_msg[9]),
    .ZN(_278_));
 OAI21_X1 _633_ (.A(_278_),
    .B1(_233_),
    .B2(_160_),
    .ZN(_279_));
 NAND2_X1 _634_ (.A1(_279_),
    .A2(_236_),
    .ZN(_280_));
 NAND2_X1 _635_ (.A1(req_msg[25]),
    .A2(req_rdy),
    .ZN(_281_));
 NAND2_X1 _636_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[9] ),
    .ZN(_282_));
 NAND3_X1 _637_ (.A1(_280_),
    .A2(_281_),
    .A3(_282_),
    .ZN(_029_));
 OAI22_X1 _638_ (.A1(_150_),
    .A2(_230_),
    .B1(_233_),
    .B2(_087_),
    .ZN(_283_));
 NAND2_X1 _639_ (.A1(_283_),
    .A2(_236_),
    .ZN(_284_));
 NAND2_X1 _640_ (.A1(req_msg[26]),
    .A2(req_rdy),
    .ZN(_285_));
 NAND2_X1 _641_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[10] ),
    .ZN(_286_));
 NAND3_X1 _642_ (.A1(_284_),
    .A2(_285_),
    .A3(_286_),
    .ZN(_030_));
 NAND2_X1 _643_ (.A1(resp_msg[11]),
    .A2(_231_),
    .ZN(_287_));
 OAI21_X1 _644_ (.A(_287_),
    .B1(_085_),
    .B2(_233_),
    .ZN(_288_));
 NAND2_X1 _645_ (.A1(_288_),
    .A2(_236_),
    .ZN(_289_));
 AND2_X1 _646_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[11] ),
    .ZN(_290_));
 AOI21_X1 _647_ (.A(_290_),
    .B1(req_msg[27]),
    .B2(req_rdy),
    .ZN(_291_));
 NAND2_X1 _648_ (.A1(_289_),
    .A2(_291_),
    .ZN(_031_));
 OAI22_X1 _649_ (.A1(_153_),
    .A2(_230_),
    .B1(_233_),
    .B2(_114_),
    .ZN(_292_));
 NAND2_X1 _650_ (.A1(_292_),
    .A2(_236_),
    .ZN(_293_));
 NAND2_X1 _651_ (.A1(req_msg[28]),
    .A2(net2),
    .ZN(_294_));
 NAND2_X1 _652_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[12] ),
    .ZN(_295_));
 NAND3_X1 _653_ (.A1(_293_),
    .A2(_294_),
    .A3(_295_),
    .ZN(_032_));
 NAND2_X1 _654_ (.A1(resp_msg[13]),
    .A2(_231_),
    .ZN(_296_));
 OAI21_X1 _655_ (.A(_296_),
    .B1(_109_),
    .B2(_233_),
    .ZN(_297_));
 NAND2_X1 _656_ (.A1(_297_),
    .A2(_236_),
    .ZN(_298_));
 AND2_X1 _657_ (.A1(_240_),
    .A2(\dpath.a_lt_b$in0[13] ),
    .ZN(_299_));
 AOI21_X1 _658_ (.A(_299_),
    .B1(req_msg[29]),
    .B2(net2),
    .ZN(_300_));
 NAND2_X1 _659_ (.A1(_298_),
    .A2(_300_),
    .ZN(_033_));
 OAI22_X1 _660_ (.A1(_156_),
    .A2(_230_),
    .B1(_233_),
    .B2(_119_),
    .ZN(_301_));
 NAND2_X1 _661_ (.A1(_301_),
    .A2(_236_),
    .ZN(_302_));
 AND2_X1 _662_ (.A1(net1),
    .A2(\dpath.a_lt_b$in0[14] ),
    .ZN(_303_));
 AOI21_X1 _663_ (.A(_303_),
    .B1(req_msg[30]),
    .B2(net2),
    .ZN(_304_));
 NAND2_X1 _664_ (.A1(_302_),
    .A2(_304_),
    .ZN(_034_));
 NAND3_X1 _665_ (.A1(_128_),
    .A2(_129_),
    .A3(_231_),
    .ZN(_305_));
 OR2_X1 _666_ (.A1(_233_),
    .A2(_125_),
    .ZN(_306_));
 NAND2_X1 _667_ (.A1(_305_),
    .A2(_306_),
    .ZN(_307_));
 NAND2_X1 _668_ (.A1(_307_),
    .A2(_236_),
    .ZN(_308_));
 AND2_X1 _669_ (.A1(net1),
    .A2(\dpath.a_lt_b$in0[15] ),
    .ZN(_309_));
 AOI21_X1 _670_ (.A(_309_),
    .B1(req_msg[31]),
    .B2(net2),
    .ZN(_310_));
 NAND2_X1 _671_ (.A1(_308_),
    .A2(_310_),
    .ZN(_035_));
 DFF_X2 _672_ (.D(_000_),
    .CK(clk),
    .Q(net2),
    .QN(_003_));
 DFF_X1 _673_ (.D(_001_),
    .CK(clk),
    .Q(\ctrl.state.out[1] ),
    .QN(_311_));
 DFF_X1 _674_ (.D(_002_),
    .CK(clk),
    .Q(\ctrl.state.out[2] ),
    .QN(_312_));
 DFF_X1 _675_ (.D(_004_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[0] ),
    .QN(_313_));
 DFF_X1 _676_ (.D(_005_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[1] ),
    .QN(_314_));
 DFF_X1 _677_ (.D(_006_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[2] ),
    .QN(_315_));
 DFF_X1 _678_ (.D(_007_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[3] ),
    .QN(_316_));
 DFF_X1 _679_ (.D(_008_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[4] ),
    .QN(_317_));
 DFF_X1 _680_ (.D(_009_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[5] ),
    .QN(_318_));
 DFF_X1 _681_ (.D(_010_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[6] ),
    .QN(_319_));
 DFF_X1 _682_ (.D(_011_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[7] ),
    .QN(_320_));
 DFF_X1 _683_ (.D(_012_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[8] ),
    .QN(_321_));
 DFF_X1 _684_ (.D(_013_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[9] ),
    .QN(_322_));
 DFF_X1 _685_ (.D(_014_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[10] ),
    .QN(_323_));
 DFF_X1 _686_ (.D(_015_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[11] ),
    .QN(_324_));
 DFF_X1 _687_ (.D(_016_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[12] ),
    .QN(_325_));
 DFF_X1 _688_ (.D(_017_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[13] ),
    .QN(_326_));
 DFF_X1 _689_ (.D(_018_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[14] ),
    .QN(_327_));
 DFF_X1 _690_ (.D(_019_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in1[15] ),
    .QN(_328_));
 DFF_X1 _691_ (.D(_020_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[0] ),
    .QN(_329_));
 DFF_X1 _692_ (.D(_021_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[1] ),
    .QN(_330_));
 DFF_X1 _693_ (.D(_022_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[2] ),
    .QN(_331_));
 DFF_X1 _694_ (.D(_023_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[3] ),
    .QN(_332_));
 DFF_X1 _695_ (.D(_024_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[4] ),
    .QN(_333_));
 DFF_X1 _696_ (.D(_025_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[5] ),
    .QN(_334_));
 DFF_X1 _697_ (.D(_026_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[6] ),
    .QN(_335_));
 DFF_X1 _698_ (.D(_027_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[7] ),
    .QN(_336_));
 DFF_X1 _699_ (.D(_028_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[8] ),
    .QN(_337_));
 DFF_X1 _700_ (.D(_029_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[9] ),
    .QN(_338_));
 DFF_X1 _701_ (.D(_030_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[10] ),
    .QN(_339_));
 DFF_X1 _702_ (.D(_031_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[11] ),
    .QN(_340_));
 DFF_X1 _703_ (.D(_032_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[12] ),
    .QN(_341_));
 DFF_X1 _704_ (.D(_033_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[13] ),
    .QN(_342_));
 DFF_X1 _705_ (.D(_034_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[14] ),
    .QN(_343_));
 DFF_X1 _706_ (.D(_035_),
    .CK(clk),
    .Q(\dpath.a_lt_b$in0[15] ),
    .QN(_344_));
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_113 ();
 BUF_X2 max_cap1 (.A(_240_),
    .Z(net1));
 BUF_X4 load_slew2 (.A(net2),
    .Z(req_rdy));
endmodule
